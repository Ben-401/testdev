use WORK.ALL;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use Std.TextIO.all;
use work.debugtools.all;

ENTITY ram32x1k IS
  PORT (
	 -- port-A is WRITE only
    clka : IN STD_LOGIC;
	 clka_en : in std_logic;
    wea : IN STD_LOGIC_vector(3 downto 0);
    addra : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
--    douta : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	 -- port-B is READ only
    clkb : IN STD_LOGIC;
	 clkb_en : in std_logic;
    addrb : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
--    dinb : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END ram32x1k;

architecture behavioural of ram32x1k is

  type ram_t is array (0 to 1023) of std_logic_vector(31 downto 0);
  signal ram : ram_t := (
    0 => x"02020202", 1 => x"03030303",
    others => x"07070707");

begin  -- behavioural

  process(clka, clka_en,
          wea, dina, addra, ram)
  begin
    if(rising_edge(Clka)) then 
 	   if (Clka_en = '1') then
        if(wea(3)='1' or wea(2)='1' or wea(1)='1' or wea(0)='1') then
          ram(to_integer(unsigned(addra))) <= dina;
        end if;
--	     douta <= ram(to_integer(unsigned(addra)));
      end if;
    end if;
  end process;

  process (clkb, clkb_en,
           addrb, ram)
  begin
    if(rising_edge(Clkb)) then 
 	   if (Clkb_en = '1') then
--        if(web='1') then
--          ram(to_integer(unsigned(addrb))) <= dinb;
--        end if;
	     doutb <= ram(to_integer(unsigned(addrb)));
      end if;
    end if;
  end process;

end behavioural;

----------------------------------------------------------------------------------
----    This file is owned and controlled by Xilinx and must be used solely     --
----    for design, simulation, implementation and creation of design files     --
----    limited to Xilinx devices or technologies. Use with non-Xilinx          --
----    devices or technologies is expressly prohibited and immediately         --
----    terminates your license.                                                --
----                                                                            --
----    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
----    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
----    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
----    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
----    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
----    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
----    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
----    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
----    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
----    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
----    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
----    PARTICULAR PURPOSE.                                                     --
----                                                                            --
----    Xilinx products are not intended for use in life support appliances,    --
----    devices, or systems.  Use in such applications are expressly            --
----    prohibited.                                                             --
----                                                                            --
----    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
----    All rights reserved.                                                    --
----------------------------------------------------------------------------------
----------------------------------------------------------------------------------
---- You must compile the wrapper file ram32x1024.vhd when simulating
---- the core, ram32x1024. When compiling the wrapper file, be sure to
---- reference the XilinxCoreLib VHDL simulation library. For detailed
---- instructions, please refer to the "CORE Generator Help".
--
---- The synthesis directives "translate_off/translate_on" specified
---- below are supported by Xilinx, Mentor Graphics and Synplicity
---- synthesis tools. Ensure they are correct for your synthesis tool(s).
--
--LIBRARY ieee;
--USE ieee.std_logic_1164.ALL;
---- synthesis translate_off
--LIBRARY XilinxCoreLib;
---- synthesis translate_on
--ENTITY ram32x1024 IS
--  PORT (
--    clka : IN STD_LOGIC;
--	 clka_en : in std_logic;
--    ena : IN STD_LOGIC;
--    wea : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
--    addra : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
--    dina : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
--    douta : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
--    clkb : IN STD_LOGIC;
--	 clkb_en : in std_logic;
--    web : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
--    addrb : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
--    dinb : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
--    doutb : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
--  );
--END ram32x1024;
--
--ARCHITECTURE ram32x1024_a OF ram32x1024 IS
---- synthesis translate_off
---- BG why syn off?
---- BG this one needs work...
--COMPONENT wrapped_ram32x1024
--  PORT (
--    clka : IN STD_LOGIC;
--    ena : IN STD_LOGIC;
--    wea : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
--    addra : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
--    dina : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
--    douta : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
--    clkb : IN STD_LOGIC;
--    web : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
--    addrb : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
--    dinb : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
--    doutb : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
--  );
--END COMPONENT;
--
---- Configuration specification
--  FOR ALL : wrapped_ram32x1024 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_3(behavioral)
--    GENERIC MAP (
--      c_addra_width => 10,
--      c_addrb_width => 10,
--      c_algorithm => 1,
--      c_axi_id_width => 4,
--      c_axi_slave_type => 0,
--      c_axi_type => 1,
--      c_byte_size => 8,
--      c_common_clk => 0,
--      c_default_data => "0",
--      c_disable_warn_bhv_coll => 0,
--      c_disable_warn_bhv_range => 0,
--      c_enable_32bit_address => 0,
--      c_family => "artix7",
--      c_has_axi_id => 0,
--      c_has_ena => 1,
--      c_has_enb => 0,
--      c_has_injecterr => 0,
--      c_has_mem_output_regs_a => 0,
--      c_has_mem_output_regs_b => 0,
--      c_has_mux_output_regs_a => 0,
--      c_has_mux_output_regs_b => 0,
--      c_has_regcea => 0,
--      c_has_regceb => 0,
--      c_has_rsta => 0,
--      c_has_rstb => 0,
--      c_has_softecc_input_regs_a => 0,
--      c_has_softecc_output_regs_b => 0,
--      c_init_file => "BlankString",
--      c_init_file_name => "ram32x1024.mif",
--      c_inita_val => "0",
--      c_initb_val => "0",
--      c_interface_type => 0,
--      c_load_init_file => 1,
--      c_mem_type => 2,
--      c_mux_pipeline_stages => 0,
--      c_prim_type => 1,
--      c_read_depth_a => 1024,
--      c_read_depth_b => 1024,
--      c_read_width_a => 32,
--      c_read_width_b => 32,
--      c_rst_priority_a => "CE",
--      c_rst_priority_b => "CE",
--      c_rst_type => "SYNC",
--      c_rstram_a => 0,
--      c_rstram_b => 0,
--      c_sim_collision_check => "ALL",
--      c_use_bram_block => 0,
--      c_use_byte_wea => 1,
--      c_use_byte_web => 1,
--      c_use_default_data => 0,
--      c_use_ecc => 0,
--      c_use_softecc => 0,
--      c_wea_width => 4,
--      c_web_width => 4,
--      c_write_depth_a => 1024,
--      c_write_depth_b => 1024,
--      c_write_mode_a => "WRITE_FIRST",
--      c_write_mode_b => "WRITE_FIRST",
--      c_write_width_a => 32,
--      c_write_width_b => 32,
--      c_xdevicefamily => "artix7"
--    );
---- synthesis translate_on
--BEGIN
---- synthesis translate_off
--U0 : wrapped_ram32x1024
--  PORT MAP (
--    clka => clka,
--    ena => ena,
--    wea => wea,
--    addra => addra,
--    dina => dina,
--    douta => douta,
--    clkb => clkb,
--    web => web,
--    addrb => addrb,
--    dinb => dinb,
--    doutb => doutb
--  );
---- synthesis translate_on
--
--END ram32x1024_a;
