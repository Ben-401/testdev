library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use work.debugtools.all;

-- this component was created with pngprepare

entity charrom is
  port (Clk : in std_logic;
        Clk_en : in std_logic;
        address : in integer range 0 to 4095;
        -- chip select, active low       
--        cs : in std_logic;
        data_o : out std_logic_vector(7 downto 0);

--        writeclk : in std_logic;
        -- Yes, we do have a write enable, because we allow modification of ROMs
        -- in the running machine, unless purposely disabled.  This gives us
        -- something like the WOM that the Amiga had.
        writecs : in std_logic;
        we : in std_logic;
        writeaddress : in unsigned(11 downto 0);
        data_i : in std_logic_vector(7 downto 0)
    );
  end charrom;

architecture Behavioral of charrom is

-- 4K x 8bit pre-initialised RAM for character ROM

type ram_t is array (0 to 4095) of std_logic_vector(7 downto 0);
signal ram : ram_t := (

-- end of upper-template
x"78",x"cc",x"dc",x"dc",x"c0",x"cc",x"7c",x"00",
-- [ ****   ]
-- [**  **  ]
-- [** ***  ]
-- [** ***  ]
-- [**      ]
-- [**  **  ]
-- [ *****  ]
-- [        ]
x"78",x"cc",x"cc",x"fc",x"cc",x"cc",x"cc",x"00",
-- [ ****   ]
-- [**  **  ]
-- [**  **  ]
-- [******  ]
-- [**  **  ]
-- [**  **  ]
-- [**  **  ]
-- [        ]
x"f8",x"cc",x"cc",x"f8",x"cc",x"cc",x"fc",x"00",
-- [*****   ]
-- [**  **  ]
-- [**  **  ]
-- [*****   ]
-- [**  **  ]
-- [**  **  ]
-- [******  ]
-- [        ]
x"78",x"cc",x"cc",x"c0",x"c0",x"cc",x"7c",x"00",
-- [ ****   ]
-- [**  **  ]
-- [**  **  ]
-- [**      ]
-- [**      ]
-- [**  **  ]
-- [ *****  ]
-- [        ]
x"f8",x"cc",x"cc",x"cc",x"cc",x"cc",x"f8",x"00",
-- [*****   ]
-- [**  **  ]
-- [**  **  ]
-- [**  **  ]
-- [**  **  ]
-- [**  **  ]
-- [*****   ]
-- [        ]
x"fc",x"cc",x"c0",x"f0",x"c0",x"cc",x"fc",x"00",
-- [******  ]
-- [**  **  ]
-- [**      ]
-- [****    ]
-- [**      ]
-- [**  **  ]
-- [******  ]
-- [        ]
x"fc",x"cc",x"c0",x"f0",x"c0",x"c0",x"c0",x"00",
-- [******  ]
-- [**  **  ]
-- [**      ]
-- [****    ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [        ]
x"7c",x"cc",x"c0",x"dc",x"cc",x"cc",x"7c",x"00",
-- [ *****  ]
-- [**  **  ]
-- [**      ]
-- [** ***  ]
-- [**  **  ]
-- [**  **  ]
-- [ *****  ]
-- [        ]
x"cc",x"cc",x"cc",x"fc",x"cc",x"cc",x"cc",x"00",
-- [**  **  ]
-- [**  **  ]
-- [**  **  ]
-- [******  ]
-- [**  **  ]
-- [**  **  ]
-- [**  **  ]
-- [        ]
x"fc",x"30",x"30",x"30",x"30",x"30",x"fc",x"00",
-- [******  ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [******  ]
-- [        ]
x"fc",x"cc",x"0c",x"0c",x"cc",x"cc",x"f8",x"00",
-- [******  ]
-- [**  **  ]
-- [    **  ]
-- [    **  ]
-- [**  **  ]
-- [**  **  ]
-- [*****   ]
-- [        ]
x"cc",x"cc",x"d8",x"f0",x"d8",x"cc",x"cc",x"00",
-- [**  **  ]
-- [**  **  ]
-- [** **   ]
-- [****    ]
-- [** **   ]
-- [**  **  ]
-- [**  **  ]
-- [        ]
x"c0",x"c0",x"c0",x"c0",x"c0",x"cc",x"fc",x"00",
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**  **  ]
-- [******  ]
-- [        ]
x"c6",x"ee",x"fe",x"fe",x"d6",x"c6",x"c6",x"00",
-- [**   ** ]
-- [*** *** ]
-- [******* ]
-- [******* ]
-- [** * ** ]
-- [**   ** ]
-- [**   ** ]
-- [        ]
x"cc",x"cc",x"ec",x"fc",x"dc",x"cc",x"cc",x"00",
-- [**  **  ]
-- [**  **  ]
-- [*** **  ]
-- [******  ]
-- [** ***  ]
-- [**  **  ]
-- [**  **  ]
-- [        ]
x"78",x"cc",x"cc",x"cc",x"cc",x"cc",x"7c",x"00",
-- [ ****   ]
-- [**  **  ]
-- [**  **  ]
-- [**  **  ]
-- [**  **  ]
-- [**  **  ]
-- [ *****  ]
-- [        ]
x"f8",x"cc",x"cc",x"fc",x"c0",x"c0",x"c0",x"00",
-- [*****   ]
-- [**  **  ]
-- [**  **  ]
-- [******  ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [        ]
x"78",x"cc",x"cc",x"cc",x"d4",x"d8",x"6c",x"00",
-- [ ****   ]
-- [**  **  ]
-- [**  **  ]
-- [**  **  ]
-- [** * *  ]
-- [** **   ]
-- [ ** **  ]
-- [        ]
x"f8",x"cc",x"cc",x"f8",x"cc",x"cc",x"cc",x"00",
-- [*****   ]
-- [**  **  ]
-- [**  **  ]
-- [*****   ]
-- [**  **  ]
-- [**  **  ]
-- [**  **  ]
-- [        ]
x"7c",x"c0",x"e0",x"78",x"1c",x"1c",x"f8",x"00",
-- [ *****  ]
-- [**      ]
-- [***     ]
-- [ ****   ]
-- [   ***  ]
-- [   ***  ]
-- [*****   ]
-- [        ]
x"fc",x"30",x"30",x"30",x"30",x"30",x"30",x"00",
-- [******  ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [        ]
x"cc",x"cc",x"cc",x"cc",x"cc",x"dc",x"78",x"00",
-- [**  **  ]
-- [**  **  ]
-- [**  **  ]
-- [**  **  ]
-- [**  **  ]
-- [** ***  ]
-- [ ****   ]
-- [        ]
x"cc",x"cc",x"cc",x"58",x"78",x"30",x"30",x"00",
-- [**  **  ]
-- [**  **  ]
-- [**  **  ]
-- [ * **   ]
-- [ ****   ]
-- [  **    ]
-- [  **    ]
-- [        ]
x"c6",x"c6",x"d6",x"fe",x"fe",x"ee",x"c6",x"00",
-- [**   ** ]
-- [**   ** ]
-- [** * ** ]
-- [******* ]
-- [******* ]
-- [*** *** ]
-- [**   ** ]
-- [        ]
x"cc",x"cc",x"78",x"30",x"78",x"cc",x"cc",x"00",
-- [**  **  ]
-- [**  **  ]
-- [ ****   ]
-- [  **    ]
-- [ ****   ]
-- [**  **  ]
-- [**  **  ]
-- [        ]
x"cc",x"cc",x"dc",x"78",x"30",x"30",x"30",x"00",
-- [**  **  ]
-- [**  **  ]
-- [** ***  ]
-- [ ****   ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [        ]
x"fc",x"cc",x"18",x"30",x"60",x"ec",x"fc",x"00",
-- [******  ]
-- [**  **  ]
-- [   **   ]
-- [  **    ]
-- [ **     ]
-- [*** **  ]
-- [******  ]
-- [        ]
x"78",x"60",x"60",x"60",x"60",x"60",x"78",x"00",
-- [ ****   ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ ****   ]
-- [        ]
x"78",x"cc",x"c0",x"f0",x"60",x"60",x"fc",x"00",
-- [ ****   ]
-- [**  **  ]
-- [**      ]
-- [****    ]
-- [ **     ]
-- [ **     ]
-- [******  ]
-- [        ]
x"78",x"18",x"18",x"18",x"18",x"18",x"78",x"00",
-- [ ****   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [ ****   ]
-- [        ]
x"10",x"38",x"7c",x"38",x"38",x"38",x"38",x"00",
-- [   *    ]
-- [  ***   ]
-- [ *****  ]
-- [  ***   ]
-- [  ***   ]
-- [  ***   ]
-- [  ***   ]
-- [        ]
x"00",x"20",x"7e",x"fe",x"7e",x"20",x"00",x"00",
-- [        ]
-- [  *     ]
-- [ ****** ]
-- [******* ]
-- [ ****** ]
-- [  *     ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"38",x"38",x"38",x"38",x"38",x"00",x"38",x"00",
-- [  ***   ]
-- [  ***   ]
-- [  ***   ]
-- [  ***   ]
-- [  ***   ]
-- [        ]
-- [  ***   ]
-- [        ]
x"6c",x"6c",x"48",x"00",x"00",x"00",x"00",x"00",
-- [ ** **  ]
-- [ ** **  ]
-- [ *  *   ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"6c",x"6c",x"fe",x"6c",x"fe",x"6c",x"6c",x"00",
-- [ ** **  ]
-- [ ** **  ]
-- [******* ]
-- [ ** **  ]
-- [******* ]
-- [ ** **  ]
-- [ ** **  ]
-- [        ]
x"30",x"fc",x"c0",x"fc",x"0c",x"fc",x"30",x"00",
-- [  **    ]
-- [******  ]
-- [**      ]
-- [******  ]
-- [    **  ]
-- [******  ]
-- [  **    ]
-- [        ]
x"c4",x"cc",x"18",x"30",x"60",x"cc",x"8c",x"00",
-- [**   *  ]
-- [**  **  ]
-- [   **   ]
-- [  **    ]
-- [ **     ]
-- [**  **  ]
-- [*   **  ]
-- [        ]
x"78",x"cc",x"cc",x"78",x"e8",x"dc",x"7c",x"00",
-- [ ****   ]
-- [**  **  ]
-- [**  **  ]
-- [ ****   ]
-- [*** *   ]
-- [** ***  ]
-- [ *****  ]
-- [        ]
x"30",x"30",x"20",x"00",x"00",x"00",x"00",x"00",
-- [  **    ]
-- [  **    ]
-- [  *     ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"38",x"60",x"60",x"60",x"60",x"60",x"38",x"00",
-- [  ***   ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [  ***   ]
-- [        ]
x"70",x"18",x"18",x"18",x"18",x"18",x"70",x"00",
-- [ ***    ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [ ***    ]
-- [        ]
x"10",x"54",x"38",x"fe",x"38",x"54",x"10",x"00",
-- [   *    ]
-- [ * * *  ]
-- [  ***   ]
-- [******* ]
-- [  ***   ]
-- [ * * *  ]
-- [   *    ]
-- [        ]
x"00",x"30",x"30",x"fc",x"30",x"30",x"00",x"00",
-- [        ]
-- [  **    ]
-- [  **    ]
-- [******  ]
-- [  **    ]
-- [  **    ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"00",x"30",x"30",x"10",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [  **    ]
-- [  **    ]
-- [   *    ]
-- [        ]
x"00",x"00",x"00",x"7c",x"00",x"00",x"00",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [ *****  ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"00",x"00",x"30",x"30",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [  **    ]
-- [  **    ]
-- [        ]
x"04",x"0c",x"18",x"30",x"60",x"c0",x"80",x"00",
-- [     *  ]
-- [    **  ]
-- [   **   ]
-- [  **    ]
-- [ **     ]
-- [**      ]
-- [*       ]
-- [        ]
x"78",x"cc",x"dc",x"fc",x"ec",x"cc",x"78",x"00",
-- [ ****   ]
-- [**  **  ]
-- [** ***  ]
-- [******  ]
-- [*** **  ]
-- [**  **  ]
-- [ ****   ]
-- [        ]
x"30",x"70",x"30",x"30",x"30",x"30",x"fc",x"00",
-- [  **    ]
-- [ ***    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [******  ]
-- [        ]
x"f8",x"cc",x"0c",x"38",x"60",x"cc",x"fc",x"00",
-- [*****   ]
-- [**  **  ]
-- [    **  ]
-- [  ***   ]
-- [ **     ]
-- [**  **  ]
-- [******  ]
-- [        ]
x"f8",x"cc",x"0c",x"18",x"0c",x"cc",x"fc",x"00",
-- [*****   ]
-- [**  **  ]
-- [    **  ]
-- [   **   ]
-- [    **  ]
-- [**  **  ]
-- [******  ]
-- [        ]
x"c0",x"c0",x"d8",x"fc",x"18",x"18",x"18",x"00",
-- [**      ]
-- [**      ]
-- [** **   ]
-- [******  ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [        ]
x"fc",x"cc",x"c0",x"f8",x"0c",x"cc",x"f8",x"00",
-- [******  ]
-- [**  **  ]
-- [**      ]
-- [*****   ]
-- [    **  ]
-- [**  **  ]
-- [*****   ]
-- [        ]
x"7c",x"cc",x"c0",x"f8",x"cc",x"cc",x"7c",x"00",
-- [ *****  ]
-- [**  **  ]
-- [**      ]
-- [*****   ]
-- [**  **  ]
-- [**  **  ]
-- [ *****  ]
-- [        ]
x"fc",x"cc",x"0c",x"3c",x"0c",x"0c",x"0c",x"00",
-- [******  ]
-- [**  **  ]
-- [    **  ]
-- [  ****  ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [        ]
x"78",x"cc",x"cc",x"78",x"cc",x"cc",x"fc",x"00",
-- [ ****   ]
-- [**  **  ]
-- [**  **  ]
-- [ ****   ]
-- [**  **  ]
-- [**  **  ]
-- [******  ]
-- [        ]
x"78",x"cc",x"cc",x"7c",x"0c",x"cc",x"f8",x"00",
-- [ ****   ]
-- [**  **  ]
-- [**  **  ]
-- [ *****  ]
-- [    **  ]
-- [**  **  ]
-- [*****   ]
-- [        ]
x"00",x"30",x"30",x"00",x"30",x"30",x"00",x"00",
-- [        ]
-- [  **    ]
-- [  **    ]
-- [        ]
-- [  **    ]
-- [  **    ]
-- [        ]
-- [        ]
x"00",x"30",x"30",x"00",x"30",x"30",x"10",x"00",
-- [        ]
-- [  **    ]
-- [  **    ]
-- [        ]
-- [  **    ]
-- [  **    ]
-- [   *    ]
-- [        ]
x"00",x"18",x"30",x"60",x"30",x"18",x"00",x"00",
-- [        ]
-- [   **   ]
-- [  **    ]
-- [ **     ]
-- [  **    ]
-- [   **   ]
-- [        ]
-- [        ]
x"00",x"00",x"7c",x"00",x"7c",x"00",x"00",x"00",
-- [        ]
-- [        ]
-- [ *****  ]
-- [        ]
-- [ *****  ]
-- [        ]
-- [        ]
-- [        ]
x"00",x"30",x"18",x"0c",x"18",x"30",x"00",x"00",
-- [        ]
-- [  **    ]
-- [   **   ]
-- [    **  ]
-- [   **   ]
-- [  **    ]
-- [        ]
-- [        ]
x"fc",x"cc",x"0c",x"18",x"30",x"00",x"30",x"00" 
-- [******  ]
-- [**  **  ]
-- [    **  ]
-- [   **   ]
-- [  **    ]
-- [        ]
-- [  **    ]
-- [        ]
,
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00" 
-- start of lower template
);

begin

--process for read and write operation.
-- BG changed some functional description
PROCESS(Clk, ram, address, Clk_en, writecs, we, data_i)

BEGIN
  data_o <= ram(address);          

  if(rising_edge(Clk)) then 
    if (Clk_en = '1') then
    if writecs='1' then
      if(we='1') then
        ram(to_integer(writeaddress)) <= data_i;
      end if;
    end if;
    end if;
  end if;
END PROCESS;

end Behavioral;
